------------------------------------------------------------------------------------------------------------------
-- 
-- File: bus_interconnect.vhd
-- 
--  ██████╗ ██╗   ██╗███████╗ 
--  ██╔══██╗██║   ██║██╔════╝ 
--  ██████╔╝██║   ██║███████╗ 
--  ██╔══██╗██║   ██║╚════██║ 
--  ██████╔╝╚██████╔╝███████║ 
--  ╚═════╝  ╚═════╝ ╚══════╝ 
-- 
-- Descrição : Interconectador de Barramento (Bus Interconnect) para o SoC RISC-V.
--             Realiza a decodificação de endereços e roteamento de dados entre 
--             o Processador (Mestre) e os componentes endereçáveis (ROM, RAM, UART).
-- 
-- Autor     : [André Maiolini]
-- Data      : [30/12/2025]    
--
------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-------------------------------------------------------------------------------------------------------------------
-- ENTIDADE: Definição da interface do Interconectador de Barramento (BUS INTERCONNECT)
-------------------------------------------------------------------------------------------------------------------

entity bus_interconnect is
    port (
        -- ========================================================================================
        -- 1. INTERFACE COM O PROCESSADOR (CORE)
        -- ========================================================================================

        -- Barramento de Instruções (IMem - Fetch)
        imem_addr_i         : in  std_logic_vector(31 downto 0);
        imem_data_o         : out std_logic_vector(31 downto 0);

        -- Barramento de Dados (DMem - Load/Store)
        dmem_addr_i         : in  std_logic_vector(31 downto 0);
        dmem_data_i         : in  std_logic_vector(31 downto 0); -- Dados para escrita
        dmem_we_i           : in  std_logic_vector( 3 downto 0); -- Write Enable
        dmem_data_o         : out std_logic_vector(31 downto 0); -- Dados lidos

        -- ========================================================================================
        -- 2. INTERFACES PARA COMPONENTES (MEMÓRIAS E PERIFÉRICOS)
        -- ========================================================================================

        -- Interface: Boot ROM (Dual Port)

        rom_addr_a_o        : out std_logic_vector(31 downto 0);
        rom_data_a_i        : in  std_logic_vector(31 downto 0);
        rom_addr_b_o        : out std_logic_vector(31 downto 0);
        rom_data_b_i        : in  std_logic_vector(31 downto 0);
        rom_sel_b_o         : out std_logic; -- Seleção para leitura de dados

        -- Interface: RAM (Dual Port)

        ram_addr_a_o        : out std_logic_vector(31 downto 0);
        ram_data_a_i        : in  std_logic_vector(31 downto 0);
        ram_addr_b_o        : out std_logic_vector(31 downto 0);
        ram_data_b_i        : in  std_logic_vector(31 downto 0); -- Leitura
        ram_data_b_o        : out std_logic_vector(31 downto 0); -- Escrita
        ram_we_b_o          : out std_logic_vector( 3 downto 0);
        ram_sel_b_o         : out std_logic;

        -- Interface: UART

        uart_addr_o         : out std_logic_vector(3 downto 0);
        uart_data_i         : in  std_logic_vector(31 downto 0);
        uart_data_o         : out std_logic_vector(31 downto 0);
        uart_we_o           : out std_logic;
        uart_sel_o          : out std_logic

    );
end entity;

-------------------------------------------------------------------------------------------------------------------
-- ENTIDADE: Definição da interface do Interconectador de Barramento (BUS INTERCONNECT)
-------------------------------------------------------------------------------------------------------------------

architecture rtl of bus_interconnect is
    -- Sinais internos de decodificação para o lado de DADOS (DMem)
    signal s_dmem_sel_rom  : std_logic;
    signal s_dmem_sel_uart : std_logic;
    signal s_dmem_sel_ram  : std_logic;

    -- Sinais internos de decodificação para o lado de INSTRUÇÕES (IMem)
    signal s_imem_sel_rom  : std_logic;
    signal s_imem_sel_ram  : std_logic;

begin

    -- -------------------------------------------------------------------------
    -- 1. DECODIFICAÇÃO DE ENDEREÇOS (Memory Map)
    -- -------------------------------------------------------------------------
    -- ROM:  0x00000000 (0x0...)
    -- UART: 0x10000000 (0x1...)
    -- RAM:  0x80000000 (0x8...)

    -- Lado de Dados
    s_dmem_sel_rom  <= '1' when dmem_addr_i(31 downto 28) = x"0" else '0';
    s_dmem_sel_uart <= '1' when dmem_addr_i(31 downto 28) = x"1" else '0';
    s_dmem_sel_ram  <= '1' when dmem_addr_i(31 downto 28) = x"8" else '0';

    -- Lado de Instruções (Baseado no bit 31 para distinguir ROM de RAM)
    s_imem_sel_rom  <= '1' when imem_addr_i(31 downto 28) = x"0" else '0';
    s_imem_sel_ram  <= '1' when imem_addr_i(31 downto 28) = x"8" else '0';

    -- -------------------------------------------------------------------------
    -- 2. ROTEAMENTO PARA COMPONENTES (Saídas)
    -- -------------------------------------------------------------------------
    -- ROM
    rom_addr_a_o <= imem_addr_i;
    rom_addr_b_o <= dmem_addr_i;
    rom_sel_b_o  <= s_dmem_sel_rom;

    -- RAM
    ram_addr_a_o <= imem_addr_i;
    ram_addr_b_o <= dmem_addr_i;
    ram_data_b_o <= dmem_data_i;
    ram_we_b_o   <= dmem_we_i when s_dmem_sel_ram = '1' else (others => '0');
    ram_sel_b_o  <= s_dmem_sel_ram;

    -- UART
    uart_addr_o  <= dmem_addr_i(3 downto 0);
    uart_data_o  <= dmem_data_i;
    uart_we_o    <= '1' when (s_dmem_sel_uart = '1' and unsigned(dmem_we_i) > 0) else '0';
    uart_sel_o   <= s_dmem_sel_uart;

    -- -------------------------------------------------------------------------
    -- 3. MULTIPLEXAÇÃO DE RETORNO AO PROCESSADOR (Leitura)
    -- -------------------------------------------------------------------------

    -- Mux de Instrução (IMem)
    -- Só retorna dado se estiver estritamente na faixa da ROM ou RAM
    imem_data_o <= rom_data_a_i when s_imem_sel_rom = '1' else 
                   ram_data_a_i when s_imem_sel_ram = '1' else 
                   (others => '0'); -- Retorna 0 para endereços inválidos (como 0x5...)

    -- Mux de Dados (DMem)
    process (s_dmem_sel_rom, s_dmem_sel_uart, s_dmem_sel_ram, 
            rom_data_b_i, uart_data_i, ram_data_b_i)
    begin
        if s_dmem_sel_rom = '1' then
            dmem_data_o <= rom_data_b_i;
        elsif s_dmem_sel_uart = '1' then
            dmem_data_o <= uart_data_i;
        elsif s_dmem_sel_ram = '1' then
            dmem_data_o <= ram_data_b_i;
        else
            dmem_data_o <= (others => '0');
        end if;
    end process;

end architecture;

------------------------------------------------------------------------------------------------------------------