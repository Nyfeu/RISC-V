------------------------------------------------------------------------------------------------------------------
--
-- File: datapath.vhd
--
--   ██████╗  █████╗ ████████╗ █████╗ ██████╗  █████╗ ████████╗██╗  ██╗
--   ██╔══██╗██╔══██╗╚══██╔══╝██╔══██╗██╔══██╗██╔══██╗╚══██╔══╝██║  ██║
--   ██║  ██║███████║   ██║   ███████║██████╔╝███████║   ██║   ███████║
--   ██║  ██║██╔══██║   ██║   ██╔══██║██╔═══╝ ██╔══██║   ██║   ██╔══██║
--   ██████╔╝██║  ██║   ██║   ██║  ██║██║     ██║  ██║   ██║   ██║  ██║
--   ╚═════╝ ╚═╝  ╚═╝   ╚═╝   ╚═╝  ╚═╝╚═╝     ╚═╝  ╚═╝   ╚═╝   ╚═╝  ╚═╝                                                             
--
-- Descrição : O Caminho de Dados (datapath) representa o 'circuito de potência' do processador RISC-V.
--             Ele contém todos os componentes estruturais responsáveis por armazenar,
--             transportar e processar os dados. Isso inclui o Contador de Programa (PC),
--             o Banco de Registradores, a Unidade Lógica e Aritmética (ALU), o Gerador
--             de Imediatos e todos os multiplexadores. Esta unidade não toma decisões;
--             ela apenas executa as operações comandadas pela Unidade de Controle.
--
-- Autor     : [André Maiolini]
-- Data      : [20/09/2025]
--
------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; 

-------------------------------------------------------------------------------------------------------------------
-- ENTIDADE: Definição da interface do Caminho de Dados (datapath)
-------------------------------------------------------------------------------------------------------------------

entity datapath is

    port (

        ----------------------------------------------------------------------------------------------------------
        -- Sinais e Interfaces de Memória
        ----------------------------------------------------------------------------------------------------------

        -- Sinais Globais (Clock e Mater-Reset)

        CLK_i       : in  std_logic;                                  -- Clock principal
        Reset_i     : in  std_logic;                                  -- Sinal de reset assíncrono

        -- Barramento de Memória de Instruções (IMEM)

        IMem_addr_o : out std_logic_vector(31 downto 0);              -- Endereço para a IMEM (saída do PC)
        IMem_data_i : in  std_logic_vector(31 downto 0);              -- Instrução lida da IMEM

        -- Barramento de Memória de Dados (DMEM)

        DMem_addr_o        : out std_logic_vector(31 downto 0);       -- Endereço para a DMEM 
        DMem_data_o        : out std_logic_vector(31 downto 0);       -- Dado a ser escrito na DMEM (de rs2)
        DMem_data_i        : in  std_logic_vector(31 downto 0);       -- Dado lido da DMEM
        DMem_writeEnable_o : out std_logic;                           -- Habilita escrita na DMEM

        ----------------------------------------------------------------------------------------------------------
        -- Interface com a Unidade de Controle
        ----------------------------------------------------------------------------------------------------------

        -- Entradas

        RegWrite_i         : in std_logic;                            -- Habilita escrita no Banco de Registradores
        ALUSrcA_i          : in std_logic_vector(1 downto 0);         -- Seleciona a 1ª fonte da ALU
        ALUSrcB_i          : in std_logic;                            -- Seleciona a 2ª fonte da ALU (Reg vs Imm)
        MemtoReg_i         : in std_logic;                            -- Seleciona a fonte de escrita no registrador (ALU vs Mem)
        MemWrite_i         : in std_logic;                            -- Habilita escrita na memória (DMEM)
        PCSrc_i            : in std_logic_vector(1 downto 0);         -- Comando para o MUX do PC
        ALUControl_i       : in std_logic_vector(3 downto 0);         -- Código de 4 bits para a operação da ALU
        WriteDataSource_i  : in std_logic;                            -- Habilita PC+4 como fonte de escrita (para JAL/JALR)

        -- Saídas

        Instruction_o  : out std_logic_vector(31 downto 0);           -- Envia a instrução para o controle
        ALU_Zero_o     : out std_logic;                               -- Envia a flag Zero para o controle
        ALU_Negative_o : out std_logic                                -- Envia a flag Negative para o controle
    
    );

end entity;

-------------------------------------------------------------------------------------------------------------------
-- ARQUITETURA: Implementação do Caminho de Dados (datapath)
-------------------------------------------------------------------------------------------------------------------

architecture rtl of datapath is

    -- ============== DECLARAÇÃO DOS SINAIS INTERNOS DO DATAPATH ==============

    signal s_pc_current           : std_logic_vector(31 downto 0) := (others => '0');     -- Contador de Programa (PC) atual
    signal s_pc_next              : std_logic_vector(31 downto 0) := (others => '0');     -- Próximo valor do PC
    signal s_pc_plus_4            : std_logic_vector(31 downto 0) := (others => '0');     -- PC + 4 (endereço da próxima instrução)
    signal s_instruction          : std_logic_vector(31 downto 0) := (others => '0');     -- Instrução lida da memória (IMEM)
    signal s_read_data_1          : std_logic_vector(31 downto 0) := (others => '0');     -- Dados lidos do primeiro registrador (rs1)
    signal s_read_data_2          : std_logic_vector(31 downto 0) := (others => '0');     -- Dados lidos do segundo registrador (rs2)
    signal s_immediate            : std_logic_vector(31 downto 0) := (others => '0');     -- Imediato estendido (32 bits)
    signal s_alu_in_a             : std_logic_vector(31 downto 0) := (others => '0');     -- Primeiro operando da ALU
    signal s_alu_in_b             : std_logic_vector(31 downto 0) := (others => '0');     -- Segundo operando da ALU (registrador ou imediato)
    signal s_alu_result           : std_logic_vector(31 downto 0) := (others => '0');     -- Resultado da ALU (32 bits)
    signal s_write_back_data      : std_logic_vector(31 downto 0) := (others => '0');     -- Dados a serem escritos de volta no banco de registradores
    signal s_load_unit_out        : std_logic_vector(31 downto 0) := (others => '0');     -- Sinal de saida da load_unit
    signal s_alu_zero             : std_logic := '0';                                     -- Flag "Zero" da ALU
    signal s_branch_or_jal_addr   : std_logic_vector(31 downto 0) := (others => '0');     -- Endereço para Branch e JAL
    signal s_alu_negative         : std_logic := '0';                                     -- Flag "Negative" da ALU
    signal s_store_unit_out       : std_logic_vector(31 downto 0) := (others => '0');     -- Dado preparado para DMEM

begin

    -- Saídas para o control path

        Instruction_o <= s_instruction;
        ALU_Zero_o    <= s_alu_zero;
        ALU_Negative_o <= s_alu_negative;

    -- ============== Estágio de Busca (FETCH) ===============================================

        -- Contador de Programa (PC) 
        -- - Registrador de 32 bits com reset assíncrono

            PC_REGISTER:process(CLK_i, Reset_i)
            begin
                if Reset_i = '1' then
                    s_pc_current <= (others => '0');
                elsif rising_edge(CLK_i) then
                    s_pc_current <= s_pc_next;
                end if;
            end process;

        -- O PC atual busca a instrução na memória (IMEM)

            IMem_addr_o <= s_pc_current;
            s_instruction <= IMem_data_i;

    -- ============== Estágio de Decodificação (DECODE) ======================================

        -- - Gerador de Imediatos (Immediate Generator)
        -- -- Extrai e estende o imediato da instrução para 32 bits

            U_IMM_GEN: entity work.imm_gen port map (
                Instruction_i => s_instruction, 
                Immediate_o => s_immediate
            );

        -- Os endereços rs1 e rs2 da instrução são enviados ao Banco de Registradores,
        -- que fornece os dados dos registradores de forma combinacional.

            U_REG_FILE: entity work.reg_file
                port map (
                    clk_i        => CLK_i,                            -- Clock do processador
                    RegWrite_i   => RegWrite_i,                       -- Habilita escrita no banco de registradores
                    ReadAddr1_i  => s_instruction(19 downto 15),      -- rs1 (bits [19:15]) - 5 bits
                    ReadAddr2_i  => s_instruction(24 downto 20),      -- rs2 (bits [24:20]) - 5 bits
                    WriteAddr_i  => s_instruction(11 downto 7),       -- rd  (bits [11: 7]) - 5 bits
                    WriteData_i  => s_write_back_data,                -- Dados a serem escritos (da ALU ou da memória) - 32 bits
                    ReadData1_o  => s_read_data_1,                    -- Dados lidos do registrador rs1 (32 bits)
                    ReadData2_o  => s_read_data_2                     -- Dados lidos do registrador rs2 (32 bits)
                );

    -- ============== Estágio de Execução (EXECUTE) ==========================================

        -- O Mux ALUSrcB seleciona a segunda entrada da ULA:
        -- Se s_alusrc_b='0' (R-Type, Branch), usa o valor do registrador s_read_data_2.
        -- Se s_alusrc_b='1' (I-Type, Load, Store), usa a constante s_immediate.
    
            s_alu_in_b <= s_read_data_2 when ALUSrcB_i = '0' else s_immediate;

            with ALUSrcA_i select
                s_alu_in_a <= s_read_data_1    when "00", -- Padrão (rs1)
                            s_pc_current     when "01",   -- AUIPC (PC)
                            x"00000000"      when "10",   -- LUI (Zero)
                            s_read_data_1    when others;

        -- A ULA executa a operação comandada pelo s_alu_control.
        -- O resultado (s_alu_result) pode ser um valor aritmético, um endereço de memória ou um resultado de comparação.

            U_ALU: entity work.alu
                port map (
                    A_i => s_alu_in_a,
                    B_i => s_alu_in_b,
                    ALUControl_i => ALUControl_i,
                    Result_o => s_alu_result,
                    Zero_o => s_alu_zero,
                    Negative_o => s_alu_negative
                );

    -- ============== Estágio de Acesso à Memória (MEMORY) ==================================

        -- Aqui ocorre o acesso à memória de dados (DMEM).
        -- Dependendo dos sinais de controle, a CPU pode ler ou escrever na memória.
                    
        -- - A ALU sempre calcula o endereço para a memória de dados.
    
            DMem_addr_o        <= s_alu_result;
    
        -- - O dado a ser escrito vem sempre de rs2.

            DMem_data_o        <= s_store_unit_out;
    
        -- - O sinal de escrita na memória vem da unidade de controle.

            DMem_writeEnable_o <= MemWrite_i;

        -- Instanciação da Unidade de Carga

            U_LOAD_UNIT: entity work.load_unit port map (
                DMem_data_i  => DMem_data_i,                          -- Palavra completa vinda da memória de dados
                Addr_LSB_i   => s_alu_result(1 downto 0),             -- 2 bits do endereço para selecionar o byte/half
                Funct3_i     => s_instruction(14 downto 12),          -- Funct3 para decodificar o tipo de load
                Data_o       => s_load_unit_out                       -- Saída de 32 bits, já tratada
            );

        -- Instanciação da Unidade de Armazenamento

            U_STORE_UNIT: entity work.store_unit port map (
                Data_from_DMEM_i => DMem_data_i,                      -- Dado já contido na memória
                WriteData_i      => s_read_data_2,                    -- Dado vem sempre de rs2
                Addr_LSB_i       => s_alu_result(1 downto 0),         -- LSBs do endereço da ALU
                Funct3_i         => s_instruction(14 downto 12),      -- Funct3 para SW/SH/SB
                Data_o           => s_store_unit_out                  -- Saída preparada para a DMEM
            );

    -- ============== Estágio de Escrita de Volta (WRITE-BACK) ===============================

        -- Mux MemtoReg: decide o que será escrito de volta no registrador
    
            s_write_back_data <= s_pc_plus_4 when WriteDataSource_i = '1' else
                s_load_unit_out when MemtoReg_i = '1' else
                s_alu_result;

    -- ============== Lógica de Cálculo do Próximo PC ======================================
    
        -- Candidato 1: Endereço sequencial (PC + 4)

            s_pc_plus_4 <= std_logic_vector(unsigned(s_pc_current) + 4);
    
        -- Candidato 2: Endereço de destino para Branch e JAL (PC + imediato)

            s_branch_or_jal_addr <= std_logic_vector(signed(s_pc_current) + signed(s_immediate));

        -- Mux final que alimenta o registrador do PC no próximo ciclo de clock
        -- - A prioridade é: Jumps têm precedência sobre Branches, que têm precedência sobre PC+4.

            with PCSrc_i select
                s_pc_next <= s_pc_plus_4           when "00", -- PC <- PC + 4
                            s_branch_or_jal_addr   when "01", -- PC <- Endereço de Branch ou JAL
                            s_alu_result           when "10", -- PC <- Endereço do JALR (rs1 + imm)
                            (others => 'X')        when others;

end architecture; -- rtl

-------------------------------------------------------------------------------------------------------------------